module RAM(input Read, input Write, input [31:0]  Data, input [8:0] Addr, output [31:0] q);

