

module neg(
	input wire [31:0] Ra,
	output wire [31:0] Rb
);

//Rb = not Ra + 1;

	
endmodule
	
